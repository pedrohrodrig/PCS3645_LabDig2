library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity sonar_fd is
    port (
        clock           : in  std_logic;
        reset           : in  std_logic;
        mensurar        : in  std_logic;
        conta_2seg      : in  std_logic;
        conta_updown    : in  std_logic;
        zera            : in  std_logic;
        zera_2seg       : in  std_logic;
        echo            : in  std_logic;
        trigger         : out std_logic;
        pwm             : out std_logic;
        saida_serial    : out std_logic;
        fim_2seg        : out std_logic;
        fim_transmissao : out std_logic
    );
end entity;

architecture sonar_fd_behavioral of sonar_fd is
    
    component trena_digital is
        port (
            clock 		      : in  std_logic;
            reset 		      : in  std_logic;
            mensurar 	      : in  std_logic;
            echo 		      : in  std_logic;
            angulo            : in  std_logic_vector(23 downto 0);
            trigger 	      : out std_logic;
            saida_serial      : out std_logic;
            pronto 		      : out std_logic;
            db_estado 	      : out std_logic_vector (6 downto 0)
        );
    end component;

    component rom_angulos_8x24 
        port (
            endereco : in  std_logic_vector(2 downto 0);
            saida    : out std_logic_vector(23 downto 0)
        ); 
    end component;

    component controle_servo is
        port (
            clock      : in  std_logic;
            reset      : in  std_logic;
            posicao    : in  std_logic_vector(2 downto 0);  
            pwm        : out std_logic;
            db_reset   : out std_logic;
            db_pwm     : out std_logic;
            db_posicao : out std_logic_vector(2 downto 0)
        );
    end component;

    component contadorg_updown_m is
        generic (
            constant M: integer := 50 -- modulo do contador
        );
        port (
            clock   : in  std_logic;
            zera_as : in  std_logic;
            zera_s  : in  std_logic;
            conta   : in  std_logic;
            Q       : out std_logic_vector (natural(ceil(log2(real(M))))-1 downto 0);
            inicio  : out std_logic;
            fim     : out std_logic;
            meio    : out std_logic 
       );
    end component;
	 
	 component contador_m is
		 generic (
			  constant M : integer := 50;  
			  constant N : integer := 6 
		 );
		 port (
			  clock : in  std_logic;
			  zera  : in  std_logic;
			  conta : in  std_logic;
			  Q     : out std_logic_vector (N-1 downto 0);
			  fim   : out std_logic
		 );
		end component;

    signal s_angulo : std_logic_vector (23 downto 0);
	 signal s_contagem_endereco : std_logic_vector (2 downto 0);

begin
    
    TRENA: trena_digital
    port map (
        clock 	          => clock,
        reset 		      => reset,
        mensurar 	      => mensurar,
        echo 		      => echo,
        angulo            => s_angulo,
        trigger 	      => trigger,
        saida_serial      => saida_serial,
        pronto 		      => fim_transmissao,
        db_estado 	      => open
    );

    ROM_ANG: rom_angulos_8x24
    port map (
        endereco => s_contagem_endereco,
        saida    => s_angulo
    );

    SERVO: controle_servo
    port map (
        clock      => clock,
        reset      => zera,
        posicao    => s_contagem_endereco,
        pwm        => pwm,
        db_reset   => open,
        db_pwm     => open,
        db_posicao => open
    );

    CONTADOR_UPDOWN: contadorg_updown_m
    generic map (
        M => 8
    )
    port map (
        clock   => clock,
        zera_as => zera,
        zera_s  => '0',
        conta   => conta_updown,
        Q       => s_contagem_endereco,
        inicio  => open,
        fim     => open,
        meio    => open
    );

    CONT_SEGUNDOS: contador_m
	generic map(
		M => 100000000, -- 2 segundos
		N => 27
	)
	port map(
		clock => clock,
		zera  => zera_2seg,
		conta => conta_2seg,
		Q     => open,
		fim   => fim_2seg  
	);
    
end architecture sonar_fd_behavioral;